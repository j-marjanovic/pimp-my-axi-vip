
package example2;

// Lorem ipsum dolor sit amet, consectetur adipiscing elit, sed do eiusmod
// tempor incididunt ut labore et dolore magna aliqua. Ut enim ad minim veniam,
// quis nostrud exercitation ullamco laboris nisi ut aliquip ex ea commodo
// consequat. Duis aute irure dolor in reprehenderit in voluptate velit esse
// cillum dolore eu fugiat nulla pariatur. Excepteur sint occaecat cupidatat non
// proident, sunt in culpa qui officia deserunt mollit anim id est laborum.

  // this function basically does nothing
  // just to test the patcher
  // add a comment in a patch
  function logic [31:0] test_function();
    logic[31:0] variable_a;
    logic[31:0] variable_b;
    int tmp;
    int tmp2;

    for (int i = 0; i < 10; i++) begin
      $display("Hello World");
    end

    // some more program

    return variable_a + variable_b;

  endfunction

endpackage;
